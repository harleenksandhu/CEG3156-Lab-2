library ieee;
use ieee.std_logic_1164.all;


library lpm;
use lpm.lpm_components.all;


entity sc_datapath is
	port(GClk, GReset: in std_logic);

end sc_datapath;


architecture rtl of sc_datapath is

end rtl;



